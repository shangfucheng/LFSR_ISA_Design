// Module Name:    ALU
// Project Name:   CSE141L
//
// Additional Comments:
//   combinational (unclocked) ALU

// includes package "Definitions"
// be sure to adjust "Definitions" to match your final set of ALU opcodes
import Definitions::*;

module ALU #(parameter W=8)(
  input        [W-1:0]   InputA,       // data inputs
                         InputB,
  input        [2:0]     OP,           // ALU opcode, part of microcode
  input                  SC_in,        // shift or carry in
  input						 parity_check,
  output logic [W-1:0]   Out,          // data output
  output logic           Zero,         // output = zero flag    !(Out)
                         Parity,       // outparity flag        ^(Out)
                         Odd,          // output odd flag        (Out[0])
//								 Neg,				// negative flag
						 SC_out        // shift or carry out
  // you may provide additional status flags, if desired
  // comment out or delete any you don't need
);

always_comb begin
// No Op = default
// add desired ALU ops, delete or comment out any you don't need
  Out = 8'b0;				                        // don't need NOOP? Out = 8'bx
  SC_out = 1'b0;		 							// 	 will flag any illegal opcodes
  if(parity_check) begin
		Out = 8'h80;
  end
  else begin
	  case(OP)
	//    ADD : {SC_out,Out} = InputA + InputB + SC_in;   // unsigned add with carry-in and carry-out
		 ADD : Out = InputA+InputB;
		 AOL : Out = {InputA[5:0],^(InputA&InputB)};	// AND ORR LSL, all in one 
	//	 AOL : Out = {InputA[7:0], SC_in};
	//    LSL : {SC_out,Out} = {InputA[7:0],SC_in};       // shift left, fill in with SC_in, fill SC_out with InputA[7]
		 BNE : Out = InputA;	// don't need out
	// for logical left shift, tie SC_in = 0
	//    RSH : {Out,SC_out} = {SC_in, InputA[7:0]};      // shift right
	//	 ORR : Out = InputA|InputB;
		 
		 XOR : Out = InputA[6:0] ^ InputB[6:0];                    // bitwise exclusive OR
	//    AND : Out = InputA & InputB;                    // bitwise AND
	//    SUB : {SC_out,Out} = InputA + (~InputB) + 1;	// InputA - InputB;
		 CMP : Out = InputA;
		 LDR : Out = InputA;
		 STR : Out = InputB;
		 
		 CLR : {SC_out,Out} = 'b0;
	  endcase
	end
end

always_comb begin
	if(parity_check) Zero = ^InputA; //~(^Out[6:0] == InputA[7]);	// using zero as parity flag, 1=error, 0 = ok
	else Zero = InputA[6:0]==InputB[6:0];	// normal zero flag

end
	
//assign Zero   = InputA==InputB;                  // reduction NOR	 Zero = !Out; 
assign Parity = ^Out;                   // reduction XOR
assign Odd    = Out[0];                 // odd/even -- just the value of the LSB
//assign Neg = SC_out;					 // negative flag

endmodule
